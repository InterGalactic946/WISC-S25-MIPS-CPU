  package Verification_tasks;

  // Task to verify that all memory locations and registers are zero post initialization.
  task VerifyPostInitialization(ref instr_memory, ref data_memory, ref regfile, ref pc, ref error);
      integer addr;
      reg [15:0] data;

      // Verify that the PC is initialized to 0x0000.
      if (pc !== expected_pc) begin
        $display("ERROR: PC not initialized to 0x0000 after reset.");
        error = 1'b1;
      end

      // Verify Data Memory (iDATA_MEM)
      for (addr = 0; addr < 65536; addr = addr + 1) begin
          data = data_memory.mem[addr]; // Accessing memory array
          if (data !== 16'h0000) begin
              $display("ERROR: Data Memory at address %0d: Expected 0x0000, Found 0x%h.", addr, data);
              error = 1'b1;
          end
      end

      // Verify Instruction Memory (iINSTR_MEM)
      for (addr = 0; addr < 65536; addr = addr + 1) begin
          data = instr_memory.mem[addr]; // Accessing memory array
          if (data !== 16'h0000) begin
              $display("ERROR: Instruction Memory at address %0d: Expected 0x0000, Found 0x%h.", addr, data);
              error = 1'b1;
          end
      end

      // Verify Register File (iRF)
      for (addr = 0; addr < 16; addr = addr + 1) begin
          // Set the source registers to each register address
          regfile.SrcReg1 = addr;
          regfile.SrcReg2 = addr;

          // Read the data from both source registers
          @(posedge clk); // wait for the next clock cycle

          if (regfile.SrcData1 !== 16'h0000) begin
              $display("ERROR: Register File Error at register %0d (SrcData1): Expected 0x0000, Found 0x%h", addr, regfile.SrcData1);
              error = 1'b1;
          end
          if (regfile.SrcData2 !== 16'h0000) begin
              $display("ERROR: Register File Error at register %0d (SrcData2): Expected 0x0000, Found 0x%h", addr, regfile.SrcData2);
              error = 1'b1;
          end
      end
  endtask

  // Task to verify the instruction fetched from the instruction memory.
  task VerifyInstructionFetched(ref expected_instr, ref actual_instr, ref mem_unit, ref instr_memory, ref expected_pc, ref pc, ref error);
      // Verify the PC.
      if (pc !== expected_pc) begin
          $display("ERROR: PC Mismatch after instruction fetch: Expected 0x%h, Found 0x%h.", expected_pc, pc);
          error = 1'b1;
      end

      // Verify the fetched instruction.
      if (actual_instr !== expected_instr) begin
          $display("ERROR: Instruction Mismatch at address 0x%h: Expected 0x%h, Found 0x%h.", pc, instr, data);
          error = 1'b1;
      end
  endtask

  // Task to verify the control signals generated by the control unit.
  task VerifyControlSignals(ref opcode, ref instr_name, )
  endtask

endpackage  