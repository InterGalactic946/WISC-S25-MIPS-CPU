`default_nettype none // Set the default as none to avoid errors

module cpu_tb();

  import Model_tasks::*;
  import Verification_tasks::*;

  ///////////////////////////
  // Stimulus of type reg //
  /////////////////////////
  logic clk, rst_n;

  ///////////////////////////////
  // Declare internal signals //
  /////////////////////////////
  logic hlt;
  logic [15:0] expected_pc;
  logic [15:0] pc;
  logic [15:0] next_pc;
  logic [15:0] instr;
  logic [3:0] opcode;
  logic [3:0] rs;
  logic [3:0] rt;
  logic [3:0] rd;
  logic [15:0] imm;
  logic [15:0] A, B;
  logic ALUSrc, MemtoReg, RegWrite, RegSrc, MemEnable, MemWrite, Branch, BR, HLT, ALUOp, Z_en, NV_en; // Control signals
  logic [15:0] reg_data;
  logic [15:0] result;
  logic [15:0] data_memory_output;
  string instr_name;
  logic [2:0] cc;            // Condition code for branch instructions
  logic [15:0] regfile [0:15];        // Register file to verify during execution
  logic [15:0] instr_memory [0:65535]; // Instruction Memory to be loaded
  logic [15:0] data_memory [0:65535]; // Data Memory to be loaded
  logic [2:0] flag_reg;               // Flag register to verify during execution
  logic Z_enable, V_enable, N_enable; // Enable flags for updating flag register
  logic Z_set, V_set, N_set;          // Flags to be set based on the result of the operation
  logic PCS;                          // Flag to determine if the next PC is the result of the ALU operation
  logic error;                        // Error flag to indicate test failure

  //////////////////////
  // Instantiate DUT //
  ////////////////////
  cpu iDUT (.clk(clk), .rst_n(rst_n), .hlt(hlt), .pc(pc));


  // Task to initialize the testbench.
  task automatic Setup();
    begin
      error = 1'b0; // Reset error flag
      regfile = '{default: 16'h0000}; // Initialize all registers to 0x0000
      
      // Initialize the PC to a starting value (e.g., 0)
      $display("Initializing CPU Testbench...");

      // Initialize all signals for the testbench.
      Initialize(.clk(clk), .rst_n(rst_n));

      // Verify that all memory locations and registers are zero post initialization.
      VerifyPostInitialization(.instr_memory(instr_memory), .data_memory(data_memory), .regfile(regfile), .pc(pc), .error(error));

      // Load instructions into memory for the CPU to execute.
      if (!error) begin
        // Load instructions into memory for the CPU to execute.
        LoadImage("instructions.img", instr_memory);

        // Load instructions into data memory for the CPU to perform memory operations.
        LoadImage("data.img", data_memory);
        
        // Print a message to indicate successful initialization.
        $display("CPU Testbench initialized successfully.");
      end else begin
        $display("ERROR: CPU Testbench initialization failed.");
        $stop();
      end
    end
  endtask

  // Test procedure to apply stimulus and check responses
  initial begin
    ///////////////////////////////
    // Initialize the testbench //
    /////////////////////////////
    Setup();

    // Run the simulation for each instruction in the instruction memory.
    repeat (instr_memory.size) begin
      @(posedge clk); // Wait for the next clock cycle

      // Fetch the current instruction from memory.
      FetchInstruction(.instr_memory(instr_memory), .pc(expected_pc), .instr(instr));

      // Verify that the instruction was fetched correctly.
      VerifyInstructionFetched(.expected_instr(instr), .actual_instr(iDUT.pc_inst), .mem_unit(iDUT.iINSTR_MEM), .instr_memory(instr_memory), .expected_pc(expected_pc), .pc(pc), .error(error));

      // Decode the instruction to extract opcode, rs, rt, rd, imm, and cc, and control signals.
      DecodeInstruction(
          .instr(instr),
          .opcode(opcode),
          .instr_name(instr_name),
          .rs(rs),
          .rt(rt),
          .rd(rd),
          .imm(imm),
          .ALUSrc(ALUSrc),
          .MemtoReg(MemtoReg),
          .RegWrite(RegWrite),
          .RegSrc(RegSrc),
          .MemEnable(MemEnable),
          .MemWrite(MemWrite),
          .Branch(Branch),
          .BR(BR),
          .HLT(HLT),
          .PCS(PCS),
          .ALUOp(ALUOp),
          .Z_en(Z_en),
          .NV_en(NV_en),
          .cc(cc)
      );

      // Verify that the control signals are correctly decoded.
      VerifyControlSignals(
        .opcode(opcode),
        .instr_name(instr_name),
        .rs(rs),
        .rt(rt),
        .rd(rd),
        .imm(imm),
        .ALUSrc(ALUSrc),
        .MemtoReg(MemtoReg),
        .RegWrite(RegWrite),
        .RegSrc(RegSrc),
        .MemEnable(MemEnable),
        .MemWrite(MemWrite),
        .Branch(Branch),
        .BR(BR),
        .HLT(HLT),
        .PCS(PCS),
        .ALUOp(ALUOp),
        .Z_en(Z_en),
        .NV_en(NV_en),
        .cc(cc),
        .control_unit(iDUT.iControlUnit),
        .error(error)
      );

      // If the HLT instruction is encountered, stop the simulation.
      if (opcode === 4'hF) begin
        $display("HLT instruction encountered. Stopping simulation.");
        $stop();
      end
      
      // Choose the correct operands for the instruction based on the opcode.
      ChooseALUOperands(
        .opcode(opcode), // Pass opcode to choose operands
        .reg_rs(rs),         // Pass source register 1
        .reg_rt(rt),         // Pass source register 2
        .reg_rd(rd),         // Pass destination register
        .imm(imm),       // Pass immediate value
        .regfile(regfile), // Pass register file
        .Input_A(A),
        .Input_B(B)
      );

      // Verify that the correct operands were chosen.
      VerifyALUOperands(
        .instr_name(instr_name), // Pass instruction
        .Input_A(A),
        .Input_B(B),
        .ALU(iDUT.iALU),
        .error(error)
      );

      // Execute the instruction based on the opcode and operands.
      ExecuteInstruction(
        .opcode(opcode), // Pass opcode to execute
        .instr_name(instr_name), // Pass instruction
        .Input_A(A), // Pass source register 1 value
        .Input_B(B), // Pass source register 2 value
        .result(result), // Pass result of the operation
        .Z_set(Z_set),
        .V_set(V_set),
        .N_set(N_set)
      );

      // Verify the result of the operation.
      VerifyExecutionResult(
        .opcode(opcode), // Pass opcode to verify result
        .instr_name(instr_name), // Pass instruction
        .Input_A(A), // Pass source register 1 value
        .Input_B(B), // Pass source register 2 value
        .result(result), // Pass result of the operation
        .Z_set(Z_set),
        .V_set(V_set),
        .N_set(N_set),
        .ALU(iDUT.iALU),
        .error(error)
      );

      // Access the memory based on the opcode and operands.
      AccessMemory(.addr(result), .data_in(regfile[rd]), .data_out(data_memory_output), .MemEnable(MemEnable), .MemWrite(MemWrite), .data_memory(data_memory));

      // Verify the memory access operation.
      VerifyMemoryAccess(
        .addr(result), // Pass address to access memory
        .instr_name(instr_name), // Pass instruction
        .data_in(regfile[rd]), // Pass data to write to memory
        .data_out(data_memory_output), // Pass data read from memory
        .mem_read(MemEnable), // Pass memory read enable signal
        .mem_write(MemWrite), // Pass memory write enable signal  
        .model_memory(data_memory), // Pass expected data memory
        .mem_unit(iDUT.iDATA_MEM),
        .error(error)
      );

      // Choose ALU_output or memory_output based on the opcode.
      reg_data = (MemtoReg) ? data_memory_output : ((PCS) ? next_pc : result);

      // Write the result back to the register file based on the opcode and operands.
      WriteBack(.regfile(regfile), .rd(rd), .input_data(reg_data), .RegWrite(RegWrite));

      // Verify the write back operation.
      VerifyWriteBack(
        .model_regfile(regfile), // Pass register file
        .instr_name(instr_name), // Pass instruction
        .reg_rd(rd), // Pass destination register
        .input_data(reg_data), // Pass data to write back
        .wr_enable(RegWrite), // Pass write enable signal
        .reg_file(iDUT.iRF),
        .error(error)
      );

      // Determine the next PC value based on the opcode and operands.
      DetermineNextPC(
        .Branch(Branch), // Pass branch flag
        .BR(BR), // Pass branch flag
        .C(cc), // Pass condition code
        .F(flag_reg), // Pass flag register
        .PC_in(expected_pc), // Pass current PC value 
        .imm(imm), // Pass immediate value
        .next_PC(next_pc),
        .Rs(reg_data) // TODO: I think this is the right net but it was missing, so double check
      );

      // Verify the next PC value.
      VerifyNextPC(
        .Branch(Branch), // Pass branch flag
        .BR(BR), // Pass branch flag
        .cc(cc), // Pass condition code
        .F(flag_reg), // Pass flag register
        .PC_in(expected_pc), // Pass current PC value
        .imm(imm), // Pass immediate value
        .next_PC(next_pc),
        .PC(iDUT.iPC),
        .error(error)
      );
    end

    // If we reached here, that means all test cases were successful
    $display("YAHOO!! All tests passed.");
    $stop();
  end

   // Expected PC value after each instruction.
  always @(posedge clk)
    if (!rst_n)
      expected_pc <= 16'h0000;
    else
      expected_pc <= next_pc;
  
  // Expected flag register at the end of each instruction.
  always @(posedge clk)
    if (!rst_n)
      flag_reg <= 3'b000;
    else if (Z_enable)
      flag_reg[2] <= Z_set;
    else if (V_enable)
      flag_reg[1] <= V_set;
    else if (N_enable)
      flag_reg[0] <= N_set;

  // Generate clock signal with 10 ns period.
  always 
    #5 clk = ~clk;

endmodule

`default_nettype wire  // Reset default behavior at the end
